module ECE_3710(input a, output b);
	assign b = a;

endmodule